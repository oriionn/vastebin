module main

import veb